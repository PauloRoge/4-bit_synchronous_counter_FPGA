library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity contador_4_bits is
    port (
        
    );
end entity contador_4_bits;

architecture hardware of contador_4_bits is
    
begin
    
    
    
end architecture hardware;